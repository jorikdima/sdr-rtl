

module selector();
	
	
	
end module